`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////////////////////////
//==================================================================================================
//  Filename      : add4.v
//  Created On    : Mon Jan  31 09:46:00 2016
//  Last Modified : 2016-02-17 08:28:17
//  Revision      : 0.1
//  Author        : Emanuel S�nchez & Ninisbeth Segovia
//  Company       : Universidad Sim�n Bol�var
//  Email         : emanuelsab@gmail.com & ninisbeth_segovia@hotmail.com
//
//  Description   : 
//==================================================================================================
////////////////////////////////////////////////////////////////////////////////////////////////////
module elbeth_add4(
    input [0:31] in,
    output [0:31] out
    );
	
	assign out = in + 4;

endmodule //elbeth_add4
